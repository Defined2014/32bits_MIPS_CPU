library verilog;
use verilog.vl_types.all;
entity ID_tb_v is
end ID_tb_v;
